.title Verification of the superposition theorem - All

vs1 1 0 dc 0
vs2 3 0 dc 2
r1 1 2 2
r2 2 4 3
r3 2 3 4

va 4 0 dc 0 ; Ammeter to measure current into R2

.end
